module mau (

    
); endmodule 