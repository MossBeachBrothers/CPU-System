module spi (); endmodule 


//Xilinx IP for SPI 

