module peripheral (); endmodule 

//Xilinx UART 



